module ex01;

initial begin
  $display(10'd001);
end

endmodule
