class Class02;

  Class01 class01 = new();

  function void method02();
    class01.method01();
  endfunction

endclass
