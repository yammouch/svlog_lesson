class Class01;

  function void method01();
    $display("Hello");
  endfunction

endclass
